vhgc
